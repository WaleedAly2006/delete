version https://git-lfs.github.com/spec/v1
oid sha256:5d83a67b82504bc01308363341bbffcf0e0615ce6ac9124664f3f448e253ca00
size 2091
