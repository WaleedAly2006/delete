version https://git-lfs.github.com/spec/v1
oid sha256:45c55f0d2a1504a19b2447823d5353410df478b2a7789062e81da82885c45cc3
size 6309
